library IEEE;
use ieee.std_logic_1164.all;
use ieee.fixed_pkg.all;

-- TEN_ARRAY is used as buffer window
-- THOUSAND_ARRAY is used as storage for testing values
package instruction_buffer_type is
type TEN_ARRAY is array (9 downto 0) of sfixed(3 downto -11);
type THOUSAND_ARRAY is array (4999 downto 0) of sfixed(3 downto -11);
end package instruction_buffer_type;

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.instruction_buffer_type.all;

entity EQ is
 port( 

        IN_FRAME : buffer TEN_ARRAY := ("000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000");
        WEIGHTS : buffer TEN_ARRAY := ("000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000","000000000000000");
        --led_low_error glows when error is less than 1%
        LED_LOW_ERROR : out std_logic ;
        CLK: in std_logic ;
        OUT_SIG : out sfixed(7 downto -22)) ;
 
end EQ;

architecture EQUALIZER of EQ is

begin
 process(CLK)
  variable EXPECTED_ARRAY : THOUSAND_ARRAY := ("100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","000100000000000","000100000000000","100100000000000","100100000000000","100100000000000","100100000000000","000100000000000","000100000000000","100100000000000","000100000000000","000100000000000");
  variable INPUT_ARRAY : THOUSAND_ARRAY := ("100011100010000","000010101000011","100100101011111","000100111010001","100100110000100","100010100100001","100111010000010","100110010110110","000001010000001","100011101001100","000100101000010","100100011010101","000100111001000","100100110011101","000100111000111","000010010111111","100000000001000","000100001100000","100100100111110","000100111110101","000010011111000","100000001001110","100011000110111","000000001101001","000011010000110","000111010101001","100000101101010","100011001111010","100111001010011","100110011111111","100110010010011","000000101001111","000011000100001","100000000110100","100011100100101","000000001011101","100011111101010","000100101101000","000010100100101","000110111110111","100000110100000","000011111110000","100100110000100","100010010111000","100111010011110","100110011001110","000000110001110","000011010001111","000111010101101","100000101010001","100011010011110","100111001100001","100110100011011","000000101010001","000011001100101","000000001100011","100011010011000","100111001001110","100110011011011","100110010000100","000000101010011","100011111111101","100010010101001","100111000011111","000000111111101","100011111111010","000100100111000","000010010011100","100000001000100","000100010011000","000010010100100","000111010010110","100000110100110","000100000111001","000010010011011","000111000001011","000110001110000","100000101111001","100011001110001","100111001110011","000000111110101","000011001111001","000000000001100","000100001100110","000010010011000","000000000101101","000100000110110","100100110101001","100010010111110","100111010110001","000000101001111","100011111111001","000100111001000","000010101110100","000111000111011","100000110001101","000011111111010","000010001001111","100000000011100","000011110001011","100100101100011","000100101100000","000010011010011","000111001000011","100000110000101","000011111011001","100100101111001","000100111001001","100100100101010","100010011011001","100111011110000","100110100000011","000000111110001","100100001000101","000100111010111","100100110010001","000100111110110","000010001001101","000111001011001","100000111100111","100010110101010","000000000110101","100011110100110","100010100010001","100111010000100","000000110000111","100011110111000","100010011011110","100111000111000","000000100010100","000011001001111","000111000110001","100000111111111","100011001000101","100111001010100","000000110011011","000011000010000","000111010101111","000110011100011","000110010111001","000110011001110","000110010111011","100001000001010","100011001111000","100000000110101","000011000100110","000111000011011","100000110111100","100011011101000","100111000100111","000000110111011","100100000000001","000100110010111","000010010011001","000000001000001","000011111110111","000010010011110","000000001010111","100011001110100","100000000100110","100100000010011","000100101100010","000010010000100","000111100001001","000110100111000","000110011100000","000110001111011","100000111010001","100011001110001","100111000110011","000000101000011","100100010010110","000100100111011","100100110000100","000100110110010","100100101111100","000100110010001","000010011011000","000111001000111","000110100000100","000110001110100","000110011101010","000110010010101","100000110101111","100011001000010","100111000100011","100110100010101","000000111101011","000011010010001","000111001100010","100000110100110","100011001110100","100111001111010","000000110011011","100011111111100","000100111001111","100100100110110","100010010101110","100111001110011","100110010100100","000000110100101","000011000100011","000000000111101","000100000010011","100100110010000","000100110111010","100100110001000","000100101011100","100100110100100","100010011010110","100111010001000","000001000000110","100100000111000","100010011101100","100000000101110","100100001001100","000100110001101","000010010111011","000111011001001","000110010111100","000110010000111","000110100110100","100000101001001","000011111110001","000010001101011","000111001001001","100000110100011","000100000010001","000010010111011","000111010000011","100000110000000","100011010110111","100111010100011","000000101101001","100100000100000","000100110000100","000010011001101","100000011000100","000011111100010","100100101001001","100010100010001","100111000101001","000000110110000","100100000000001","000100110100101","000010001100111","000111001100000","000110100110100","100000110010011","100011001100011","100000000101111","100100000000001","100010010111101","100111001001010","100110011100100","000000110001010","000011011101001","100000010010010","000100010010000","100100110000011","000100111011010","100101000000101","100010011110011","100000000010010","000011010000001","000110111111010","100000101111011","000011110110001","000010011010001","000000000101010","000100000010101","100100101010011","000100111011010","100100111000011","100010010111100","100111010100011","000000101000011","000011010100010","000000000000000","000011111111100","100100101011110","100010010100110","000000000010110","000011010110111","000111010100010","000110011011100","100000111000110","100011010010000","000000001001101","000010111111110","000111001100100","100001000010111","100011000100100","000000000110111","000011001100110","000111001100001","100001000111010","000100000100101","100101000100111","000100100000011","100100110010100","100010100001010","000000000011010","100011111010100","000100111010001","000010010100000","000000000011101","000100000000110","100100101100100","100010010101010","100111000101100","100110011010101","100110011010110","100110010001011","000000100010000","100100000100000","100010100011111","100000000011000","000011010010000","000000000110101","000011110111110","100100110111000","100010011000011","100000000010010","100011111101100","100010010110010","100000000111100","000011001011010","100000010001010","100011000011100","100000000101000","000011000011000","100000000010000","000011110100011","000010011001011","100000000100100","100010111011001","000000001001001","100100010100001","000100110110110","100100111110100","000100110001001","100100110001110","000100111001010","100100110101011","100010001100110","100111010000101","100110010110111","100110010100001","000000110011111","000011010011111","000111001111011","100000111001100","100011011011011","000000001111000","000011000111111","000111001101101","000110011110001","100000110010010","100011010100000","100111010000100","000000110010001","000011011000110","000111000101110","100000101100110","100011001010010","100000000001111","000011000100001","000111001010011","100000110011111","000011110100000","100100110001101","100010100000010","100111001101100","100110010110111","000000101011111","000011001010011","000000000010110","100011011011101","100111000100011","000001000110110","000011010100100","100000000010100","000100000011011","000010010001001","000111011100000","100000101011100","100011000110011","100000000111000","100011111101011","000100101110101","100100110101101","000100101110100","100100111011100","000100101011110","100100110100111","000100100101011","100100101110010","000100110010001","100100101101100","000100110101011","000010011101100","100000001100000","000011110111101","100100110110110","100010011000101","000000001001001","000011001010011","000111010111000","000110011101011","000110100011000","100000110010001","000011111010101","100100111111001","100010011000010","100111000110001","100110011011111","000000101110110","100100000010011","000100101010010","100100110111001","000100110001101","000010011001111","100000000000100","100011000111110","000000000000111","000011011011011","000111001111010","100000100100100","000011111010001","000010011101110","100000000010000","000100000100110","000010011110011","000110111011000","000110001110110","000110001101111","000110011100110","000110100101100","100000110101110","000100000110100","100100101110110","100010100010000","000000000011001","100100000110000","100010001101010","100111001101000","100110001100010","100110011101000","100110010100110","000000110010101","000010111100011","100000000111111","000100000100111","100100110011101","000100101010001","000010010100100","000000000010000","100011010100110","000000000111111","000011000111100","000000001110101","100011010101100","100111001011001","100110100101111","000000101101010","000011000111111","000000000011001","000100000111101","000010011100000","100000000011000","000100000110100","100100101100101","100010011000101","100111001000001","000000110110100","100100000111111","000100111001010","100100111000100","000100101110010","000010011011000","100000000010011","100011001101110","000000000100110","100011110111100","100010011011001","100111001010001","100110011011100","100110010111101","000000110110110","000011000111110","000111001111000","100000101110010","100011001100000","100110111110110","100110011110100","100110011111100","100110100111110","000000111010100","100011111000111","000100110010100","100100101011111","000100110100101","100100110000110","100010011000101","000000000011100","000011001101100","000111100011010","100000111100101","100011011011110","100111010110000","000000101010010","100100000011100","100010011010111","100111001110100","100110010101001","100110010110011","000000111001010","000011011011001","000000001001111","100011010111001","100000010010110","000011010100000","000110111101111","000110011010001","100000110010111","000100010010000","100100110011110","100010011101101","100111001010111","100110010111100","100110011001000","000000101110010","000011000010111","000111001111010","100000111110000","000011110111101","000010100100011","000111001001011","000110011000011","100000101011111","100011001111001","100111000100011","100110011100011","000000111011011","100011111010111","000100110001011","000010010010100","100000001000011","000011111101110","000010010110000","100000000011010","000100000111111","000010010111001","000000001001010","100011010001000","000000000111110","100100000100001","100010011000001","000000000111110","000011001001011","100000000011100","000100010000001","000010100001010","100000000011011","000100000101010","100100110110000","100010010011111","000000001011011","100100001100111","100010010001010","100111000000111","100110011001001","100110001011011","000000110100011","000011000010110","100000010001110","100011001111011","100111000111000","000000110101110","100011111100101","000100101110100","100100110010000","100010100110110","100000000110001","000011000110001","000000000100001","000011111111111","000010010000001","000111001100101","000110010100000","000110010100001","000110100000100","100000110010010","100011001001100","000000000111001","100011111110100","000100110111101","000010011111001","000000001001011","000100000011110","000010100101000","000000000000001","100011001101001","000000001101110","100100000100001","000100110011001","000010100001000","000000000001001","100011000001011","100111000100011","000000110101100","000011000110100","000000000100100","000011110100110","000010011011100","000111010011010","000110011011010","100000101100000","000100010000100","100100101011101","000100110101010","000010011110110","000111010000001","100000111101110","100011010000001","000000001001111","000011001100011","000111010001100","100000111011010","000100000000100","100100101110010","000100101000001","000010011100011","100000000001011","100011010100011","100000000000010","100100001111010","100010101010110","100000001001100","000011000100110","100000001001011","000011110010000","000010011011111","000110111111111","100000110010010","000100000110010","100100110011001","100010011000110","100000000011000","100100001100000","000100110010110","100100101011011","000101000001010","000010010110000","000110111111101","000110011010111","100000110000001","100011001110101","100000001001010","000011011101001","100000010011000","100011010000111","100111010111011","000000101110000","000011001111010","000000000001000","000011111010001","100100101100111","000100111000001","100100101101111","100010011101000","100111000100010","000000111000100","100011101011101","000100111011110","000010100010111","000111001101001","000110001111001","100000110110001","100011010010111","100000000100100","000011010001010","100000000100100","000011111000110","000010010110010","100000000001010","000100000011010","100100111010111","000100110101110","000010011010001","000111010111100","100000110100111","000011111110111","000010010000000","100000001011001","100011001010010","100111001110110","000000110111010","100100000111001","000101000010101","000010011010100","000000001000011","000011111110001","000010011000010","000111010010011","000110011110000","100000111100010","000011110011100","000010010000101","000111000001010","000110011010000","000110010110010","000110010110100","100000111110001","000100000110010","100100101111101","100010011010010","100111000100100","100110100000101","100110010110001","000000110110000","000011001111101","100000000101111","000100000010101","100100110111010","000100101011111","000010001111110","000111010101001","100000111010000","000011111110100","000010001111110","000111001010011","000101111111011","000110010000110","100000111110101","000011110111110","100100110100111","100010011100001","100110111101000","100110011110001","100110011011100","100110100110010","000000101111010","000011000001111","000111001101000","000110100000100","100000101111111","000011111010010","100101000000011","000100111111000","000010101010001","000000000000111","000011110111111","000010100011010","000111001000000","100000110111000","100011000101100","100111011000000","000000100011010","100011111100100","100010010110010","000000000000110","000011010000110","000111010101100","100000101011010","100011010001011","100111000110001","000000110100100","100100000100000","000100101001100","000010011110110","100000000010110","100011001100011","100000000110011","100100001100100","000100110100100","100100110011101","000100111100111","100100101100101","000100111011101","100100111001010","100010100001001","100111010111000","000000110111001","100011101001011","000100111001000","100100111001011","100010010010110","100111010101111","100110100101001","000000111001000","000011000110100","000111001111010","000110100100111","000110011100110","100000101011101","100011011001110","000000000101010","100011101110101","000100110111100","100100111111101","000100110001100","000010010101100","000000000011000","100011001001011","000000000011010","100100000010111","000100101110010","100100110111111","100010010010101","100111011011110","000000110001100","000011001110111","100000000101010","100011001000111","100111001101011","000000101011100","100011111110101","000100110001000","100100110110100","000100101101011","100100110010101","100010101000100","100111010000000","000000101110110","000011000101011","000111010010000","000110010011101","000110011101111","100000101011010","000011111110101","000010011011110","000111010001111","100000110011110","000100000100011","100100111101011","100010010000100","100000001000000","000010111101111","000111011000000","000110011001000","000110011101001","000110010110101","000110010001010","100001001100000","100011000111101","100111001111000","000000110001100","100011111100101","000100100111101","100100111001000","000100111100011","100100101110010","100010100011111","100111011110101","100110011110001","100110010111110","000000111010110","100011111111001","000100101010000","000010011100000","100000001001011","100011010100100","100111010010000","100110100011100","000000110001000","100100000111010","000100110000111","100100110110111","100010011100111","100000000100000","100011110110000","000100111000001","100100110010101","100010100101011","100111011001111","100110101001100","100110000100100","000000111011000","100011111101111","000100101011010","100100111100011","000100110111101","000010100110010","000110111111000","000110010101111","100000110011111","100011011100111","100111000101111","000000101111110","000011011100010","000111001001101","000110011100111","000110010000010","000110010100100","000110010000001","000110011100110","000110100100001","000110010100110","000110011101001","100000110111010","000100000000110","000010100011010","000111001101110","000110010001001","100000111010001","100011001110001","100000000001100","000011000101110","000000000001011","000100001010010","000010010111100","100000000001101","000011101110001","100100111001011","100010100100111","100000000011001","100011111011101","000100111111100","100100100100101","100010011010100","100111001111011","000000111001110","100011111100000","000100111001011","100100101100111","000100100111001","100100101110110","000100110010011","100100111001010","000100101101100","000010100011111","100000000110100","100011010110110","000000000001101","100011101111101","000100110011011","100100110000101","100010100001001","100110111111001","000000110100001","000011010001000","100000000111101","000100000110111","100100110000000","000100101001110","000010011001111","100000000011101","100011001011111","100000000010000","000011001011010","100000001000010","000011111101011","000010011111110","000111011010111","000110010000001","100000011111111","000100001100010","100100110001110","100010011100000","100111010010011","100110010010110","000000101101100","000011001001000","000000000111001","100011001001010","100111000101100","000000110111010","100100000011001","100010011101110","100111000110010","000000101101110","000011010110011","000000000110011","000100000010010","000010011001101","000111001111110","100000010110101","000011111111000","100100111111110","100010001010000","100111000111110","000000101101111","100011101010110","100010010101001","100111001010011","000000101100111","100100001000100","000100100100111","100100110110100","000100101010101","000010011110110","000111001010001","100000100100111","000100001100001","100100110001110","000100110000111","000010100010111","000111000011100","100000101101101","000011111010100","100100110110011","100010011111000","100111001000001","100110011111111","100110100010001","100110010101000","100110011101000","100110010110101","100110011100011","000000110101011","100100010100110","000100110110111","000010101000100","000000001000011","100011000101011","100111001110101","100110011000001","100110010111100","100110011000110","100110100000010","000000110000010","000011001011011","000111001000111","000110100000010","000110101110001","000110001110111","000110011010101","100000111110111","000100001010100","100100100111110","000100100101101","000010101001010","100000001000110","100011001010111","100111000011111","000000110100011","000011011111011","000000010110010","100011001011101","100000001111011","100100000010111","100010100000011","100000000110001","000011000011101","000000000000101","000100010001000","100100111000111","100010011011110","100111000011010","100110001111110","000000110111001","000011010101000","000000000111000","100011001111111","100111001001010","000000110000110","100100000111010","000100111000010","000010011010001","100000000001100","000100000010010","000010100001100","000000000011001","000100000001100","000010011011110","000000000000011","000011111001101","000010011111111","000000001011011","100011010001000","100110111101001","100110011011000","000000110001001","000011000101100","100000000110011","100011010100100","100111001001111","100110001100101","100110010101010","100110010010101","000000111110000","100100010100001","000100110001110","100100110000010","000100111001000","000010001111000","000111000100101","100000101100110","100011001101101","000000000100011","000011000101000","100000001101001","100011000110101","000000001001101","100011110010110","100010100110000","100000001010110","000011000000110","000111001100011","100000111000001","000100001010101","100100111110111","000100100101000","000010011011010","000111010110011","000110010011000","100000111101011","100011001110000","100000001101001","000011001100111","000111010011100","000110011011010","000110001010001","000110010101010","100000110101101","000100001110101","000010100001000","100000000000011","000100001010100","000010010001001","000111001001111","100000100111110","100011000000101","100111000110111","100110010101101","100110011110010","100110010011100","100110100000010","100110010100111","100110010111010","000000111100011","000011001001010","000000000101001","100011000110011","100000000111010","000011001110000","000111011001101","100000110010010","100011001111010","000000000011101","000011001010100","000000000011100","100011001101111","100000000000001","100011111100010","000100111110001","000010011101010","000000001101010","100011011101001","100000000011101","000011001110101","100000000110110","000011110101101","000010011110100","000111010001110","100000110000110","100011001001100","100000000111000","000011001000110","100000000000110","000011111010011","000010011100010","000111011111111","000110010101101","100000101101111","000011110111101","100100101000010","100010100001011","100111001011000","100110011110100","000000110111010","000011001100111","000111001100011","000110110001011","000110010100011","000110011001001","100000011101011","100011010110000","100111001000010","100110100010010","100110010001010","100110010110111","000000111000011","100100000010010","100010010111100","100111000000111","000000100000110","000010111111100","000000000011010","100011010010000","100000000010011","100100001100000","100010100000111","100111010000000","000000101101010","100100000111000","000100101111110","100100111010110","100010001110101","100000001000000","000011011011100","100000000011000","000011110100001","100100111000001","000100111010110","000010100010001","000111001110000","000110011011111","100000101110000","100011011000100","100111010001100","100110101000011","000000101111100","000011010100011","000111010010100","000110101100000","100000110001110","000011101110100","100100100101100","100010001111001","100111010001100","000000110101000","100011111001101","000100110110010","100100101101100","000100110010010","000010011001010","000111001101100","000110010011001","100000100111101","100011001100101","000000000101100","100100000110111","000100101010011","000010011000110","000111001010110","000110100011010","100000101110010","100011001000011","100111011000011","000000101011010","000011001110011","000111001001111","100000101000110","100011000001111","100000000100101","100011111000111","000100111110011","000010011100001","000111011001111","100000101010100","100011001011000","100111000101101","100110011000000","100110011100111","000000110110000","000011001101000","000111001001110","000110100111111","100000110001011","100010110110101","100000000010011","000011010001010","000000001100110","000100010110000","000010011100000","000111000110011","100000101100101","000011110101010","100100110101011","100010010111011","000000001100000","000011011000011","100000000000001","100011000101010","100000000010100","100011111010101","100010001010000","000000000001010","000011001010010","100000000100000","100011000110111","100111000001111","100110001000011","000000110011101","000011001110000","000111000111101","100000100110001","000011111111011","100100110111000","000101000100111","100100101100101","000100111000111","100100111011010","000100110110101","100100101110111","100010100010011","100111001110101","100110011100111","000000110111011","000011000100101","000111010101100","100000100100110","100011001111010","100000000000000","100011111011111","000100111100111","100100101110111","100010010110011","100000000011111","000011001010111","000000000100111","000100001101100","100100101110100","100010100011010","000000000011100","100100000000101","100010011011100","100000000001110","100100000111000","000100110000100","000010010011001","000111001001110","100000110010010","000100000001011","100100110100111","100010011010110","100111001100100","100110010101111","100110001111001","000000111000001","000011001010011","000111010001101","100000110101001","000011110001100","000010000110100","000110111110111","100000110101000","100011010001110","100111010010101","100110011001010","100110011110111","100110011110101","100110010100101","100110010011010","100110000101110","100110010111001","100110011001001","100110011110001","000000110001100","100100000000011","000100100100111","100100110101010","000100111001010","100100110111110","100010010101100","000000001000000","000011010101100","000111010011000","100001000101011","000011111011011","100100101011111","000100110110011","000010011001101","000111010000010","000110100010101","000110011010110","100000111001010","000011111110100","000010010111111","000000000111010","000100000011010","000010011110000","000111001101111","100000110110001","000100000000011","100100110001011","100010100100111","100111001011010","000000111010101","000011001011111","000000001100101","100011001000010","100000000011011","100100000001001","100010011011110","100111001010110","100110010011011","100110011011111","100110010101111","000001000001011","100011111000011","000100111001111","000010010011000","100000000100010","000100000001111","100100110100000","000100100110000","100100111111011","000100111011100","100100111001010","100010001000110","100111011110110","100110010101111","100110011001100","000000101101000","100011111100101","100010100000000","000000000110111","100011111111011","100010100110110","100111100000011","100110011011111","100110010000010","000000110100101","100011111111100","100010010100000","100000001011010","100011110100011","100010100000110","100111001100011","000000110000010","100011111110110","100010101001010","100111000000011","000000110111100","000011011101000","000000001011011","100011001100101","100111010100011","100110100111101","000000110011010","000011001110100","000111010101010","100000111010111","000100000110011","000010011010001","000111000110100","100000101100111","100011001010101","100000000001111","100011110000110","000100111000001","100100110100000","000100110101011","000010011010010","000000000001011","000100000011101","100100111000000","100010100000000","000000000010111","100011110000101","100010011100000","100111010100111","100110011011100","100110011101100","000000110000100","000011010000101","000111001011101","100000111000000","100011010000011","100000001010101","100100000110111","100010100101000","100000000100001","100100001000110","100010011111010","100000000010011","100100001001101","100010011001110","100111001010000","000000101011011","000011010101110","000110111111111","000110010110011","000110001101100","000110010110110","000110001110111","000110010100111","000110010011100","000110010000000","000110001000111","100000101110101","000100010000001","000010101011100","000111001000110","100000110011100","100011010000100","100111001100001","100110100001000","000000100011101","000011001100100","100000001001111","000011110000100","100100011111111","000100110001010","000010011100110","000111010110011","000110001011111","000110011100111","000110011101101","000110011010010","000110011010111","000110010101010","000110011111011","000110010010101","000110010011001","000110011111011","100000100101100","100011001111111","100000000100000","100011111100101","100010010000111","000000000111110","100011111101110","000100101110000","100100101110000","000100110010100","000010100100101","100000001011011","000100000001001","100100101000110","100010011101100","100111010001110","100110100001001","100110011011110","100110011011001","000000110100010","000011000101101","000000000000101","000011111011000","100100110110001","100010100000011","100000000010010","000011101001101","000000011011100","100011000011100","100111000110011","100110100011111","000000101110011","000011000111110","000000000100010","100011001000111","000000000000111","000011001010000","000111000101010","000110011001101","000110100010110","000110011101000","000110011011000","100000101101111","100011001000000","100111011001111","000000110011010","100100000011011","100010101010000","100111010111100","000000110000100","100011111001010","000100110001010","100100110001000","100010100000110","100111011110010","000000110011111","100100000111101","100010010000000","000000001110000","000011001001110","000111010110011","100000101011011","100011011000010","100000000000010","100011111101111","100010010101010","000000000101011","100011111010100","100010010100000","100000000010100","100011111100111","100010101011110","100000001001011","000011010110100","000111000111011","000110011100010","000110100101110","000110010010011","100000111010111","100011010000110","100111001001001","100110011011010","100110100001100","000000100110011","000011001001110","100000000001110","100011010001001","100111001110111","100110100010011","100110010101001","100110101011001","000000110100010","100011111010100","000100101100010","000010011001001","000000000010010","100011010001110","100000000000000","100011111100101","100010100001001","000000000110110","000011010101101","000000000010100","000100000000000","000010010000001","000111010000110","100000111101000","100010111111111","000000000100010","100011111101110","100010011100110","100111011110011","000000101001100","100011111101000","100010000110000","000000000101111","100011111101011","100010011101111","000000000000111","000011010100100","000111001010101","000110101000111","000110001111101","000110010110100","000110011010000","000110001001110","100000101110100","000100000000101","100100110010100","100010010011001","100111000100010","100110010011000","000000101111011","000011001100011","000111001111101","000110001111011","100000111011100","100011010000010","100111001100001","000001000001101","000011010011010","000111001001001","100000111000010","100011000000011","000000010110001","100011111110101","000100101111010","000010001110001","000000000111111","000100000010010","100100101001110","000100101011110","100100110001010","100010011110111","000000001010010","000011001000010","000111001100000","100000110110000","100011000100110","000000000011011","000011000100101","100000000101000","000011110111100","100100101111000","100010010110111","100111011010000","000000100011110","000011001100011","000111010010011","100000110001110","100011011001010","100000001100100","100011111000111","100010011010110","100111001111111","100110001110111","100110100000000","000000110100010","000011010000001","000111010011011","100000111010000","000100000010111","000010101111110","100000001100001","000100000011100","100100110101000","000100101100100","000010010010110","000111010000110","100000100000011","000011111001100","100100101110110","100010011110001","100110111100110","100110010101001","100110011010101","000000111000001","000011001100110","000000001000111","000011111110011","000010010000100","000000000001111","000100001100101","100100111100111","100010011011100","100111000100101","100110101001001","000000111000010","100011111001111","100010010111110","100000000110001","000011001100101","000111001101100","100000101011101","000100000101010","000010010110110","000000001101000","100011001101001","100111010011011","100110011101001","100110010010101","100110011000000","000000111010011","100011111111011","100010000101011","100111011010010","100110011100111","000000110010100","100011111111010","000100111110111","000010011011011","100000000000111","100011001100001","100111000110101","100110011111001","000000110110110","100100001100101","100010011010001","100111010100011","100110011110111","000000110101011","100100001001000","100010100001100","100000001100010","100100010010000","100010011010110","000000001001011","100100000001011","000100110001010","000010010001001","000000001100110","000011111101111","100100101000101","000100110110001","100100110101010","000100111011111","100100101011001","000100110010010","000010100100000","000111011011001","000110011001000","100000110101010","000100000011010","000010011100011","000000000110100","100011001110110","000000000101110","000011010101010","000000000001011","100011001011100","100111010110111","000000101001101","000011000000111","100000001010000","000011111110101","100101000000010","000101000101011","100100101101001","100010101010010","100000001001010","100100000000110","000100100101010","000010010101111","000111010101101","000110011000010","000110011001000","100000111011010","100011010001010","100111010111101","100110010110101","000000101111100","000011010011001","000000001010000","100011000100000","100000000000010","100100000100000","000100101001010","100100110010001","000100111010111","100100110101111","000100110001110","000010011110100","000111010011110","100000111110101","000100000001100","100100110001100","000100110001111","100100101011111","100010011100100","100000000110101","100011111101110","100010010101111","100000000001110","000011010011001","000111000000100","000110010000111","100001001100000","000100000100001","000010010001100","100000000010000","100011000100101","100111001100011","000000101111101","000011000101111","000111001010110","000110011110011","000110001101010","000110011001000","000110011111111","000110001110000","100000101101110","100011000111010","100000000111001","000011000000100","000000000011100","100011000110010","000000000100101","100011111001110","100010100011001","000000000100101","100100000100101","100010011110001","100000001100100","100011110111000","100010011000001","100111000100101","000000111111011","000011000011100","000000000101001","100011001100111","100111000101011","000000111100001","100011111001010","000100101100100","100100110100001","000100110101010","100100011001101","100010001111101","100110111010000","100110010110001","000000110100111","100011111011000","000100101110111","100100101001001","000100110001111","000010001110011","000111010011110","000110001100111","100001000010001","000100000010010","000010010001111","100000000111010","000011111110101","000010010101101","000111001010111","100000110000111","100011010110010","100000001001111","100100010000111","100010011100110","000000000101011","100100000101101","000100110111010","000010011101111","000111010100110","100000101011001","000011111010011","100100111010001","100010011001001","100000000101011","000011011000100","000000001011001","000100000000110","100100110110101","000100110111010","000010010100010","100000000001000","000011111011101","100100110010010","100010010000011","000000000110000","100011110110101","000100101011110","000010011011000","100000000111111","100011001001101","000000000010101","000011010111010","000111010101101","000110011110111","100000110111010","100011010000101","100000010000100","100100000011101","000100100110101","000010100001001","000111010100000","000110011010101","100000110110010","000100000001001","000010100110100","000111010111101","100000110110110","000100000001010","100100111100010","000100110110011","100100101101001","100010010010010","100111011001001","100110010101100","000000101100001","100100000011000","000100111001100","100100110000110","000100110001110","100100101110010","100010001100010","100111010001110","000000101000010","000011000011011","000111000101001","000110010100001","000110011110010","000110001000101","000110011011100","100000111001100","100011000011111","100111010011101","100110011001100","100110100001001","100110011111000","000000110001000","100100000001110","000100101110111","100100101010000","000100110111101","000010101000100","000111001010100","000110100010001","000110001000100","000110011110110","100000110000001","000011111100111","100100101101100","000100111010010","100100101010110","000100110110100","100100101110010","000100101101101","000010010000101","100000000010001","100011001011010","000000000111101","000011000110011","100000000011111","000100011000000","100100111000001","000101000010101","100100101011011","100010011110000","100111001101101","000000110001011","100011111100001","000100111110010","000010001100010","000111011101001","000110011111111","100000110111101","100011001101110","100111001010010","100110010111001","000000111100111","000011010101101","000111001001111","100000110100010","100011000110110","000000000000111","000011010101111","000111000111001","000110011101011","000110011011111","000110100100110","100000111110000","000100000000000","100100110010110","100010101100100","100111000010101","000001001001111","100100000001111","100010010111010","100111010000100","100110010110011","000000110000001","100100000000110","000101000000010","100100111010000","100010011110010","100111001101011","100110011010101","100110001101111","100110001001001","000000101011010","100100000101001","000100110111011","100100110110010","100010001001011","000000001101001","000011010001010","000000000100100","100011001111100","100111000110100","100110010000011","000000110100010","000011011100011","000000000101011","000011111111000","000010011100100","000111010101101","100000110110011","100011001101011","000000010011001","100100000011110","000100111010110","100100101100100","100010001100101","100111001000100","000000011111001","100100000110111","100010010101011","000000000010000","100011110000000","100010001110001","000000000100000","100011111111010","000100100110101","000010101000101","000000000001000","100011011001010","000000000011100","000011001101101","100000000100100","000100000011111","100100111000111","100010100100100","100111011011000","100110011100100","100110011110101","100110010110000","000000100111000","100100000001101","100010100101110","000000001110101","100100000000111","100010001111101","000000000100000","000011010100001","000111000011011","100000101001000","100011000001000","100000010000110","100100000001011","100010011110111","000000000001010","100100000110111","000100110101011","100100101110010","100010010111100","100000000000111","000011000010010","000000000000011","100011010001000","100000001010010","000011001100010","000111001011000","100000110001101","100011000100110","000000000100101","100011110101011","100010011111100","100111010011110","100110011010010","000000111110011","000011010111010","000111001011110","000110010100110","100000111111100","000100000101011","100100110011000","100010100011001","100000000010101","000010111101111","000000000011011","100011001110001","000000001101001","100100001011000","000100111011000","000010011010110","000000000000101","100011000110111","100111000011001","000000101010100","000011010111011","100000001001110","000011110111010","000010010100001","000111010010110","000110010000111","100000110000011","100011001001011","100111001011100","000000110111101","100100001001011","100010010001011","000000000000111","000011010010101","000111000100110","100000110010110","100011000101101","000000001000001","100100000000101","000100100100001","000010010000101","000000000001110","000100000110011","100100101111011","100010011110100","000000010010001","100011111111011","000100111010001","100100110110100","000100101010001","000010011111001","000000001000011","000100001110110","100100110111011","000100100110000","100100100110000","100010010111011","100111010101111","000000101110101","000011000110010","000111010110001","100000101110011","000100000001111","100100110001010","100010100000010","100111000100110","100110010110110","000000110001000","100100000001011","100010011010011","100000000111001","000011010010110","000000001011010","100010111000110","100111001000101","000000101100100","000011001110011","000111000100101","100000111000001","000011111010101","000010010010110","000000000011000","100011010101110","000000000101011","000011010011001","000111010101001","000110011001011","100000101110001","000100001110100","100100110010110","000100110001110","000010100111111","100000010100010","000011111100010","000010101101010","000111001000111","100000110111101","100011010110101","000000000110011","100100010001000","100010100000000","000000000100100","100100000000000","000100111000010","000010011010100","000111010010010","100000111101100","100011001011000","100111011001011","100110010011010","000000110000101","100011111010101","100010011101111","100111001010001","100110010001000","100110101001101","100110101000101","000000100100010","000011010011101","000111010000000","000110010011111","100000100111000","100011001011101","100000001100110","100100001000010","000100100111111","100100101011011","100010011110011","100111010110010","000000101110100","100100000110110","100010010010101","100111001000111","100110010111001","100110010110001","100110011001010","000000101011100","000011010001001","100000000110101","100011010101011","100000001000101","000011010011110","000000000111111","100011011011000","100111001101111","100110010111100","000000101110010","000011010010111","000111001110110","100000110100011","100011010001010","000000000101011","000011010011101","000111010000100","100000110101001","100011000101010","100000000111010","000011001101111","000111011000000","000110011000000","100000111010000","000100001111101","100100110101001","100010010110000","100000000110100","100011111101101","100010010101110","100111001100110","100110010110111","100110001111110","100110100100111","000000110100110","100100010000000","100010011001010","000000001111101","000011010100011","000111001100101","100000110101111","100011001000100","000000001000100","100011111111111","100010001100100","100000000110100","000010111100101","000111000110101","000110010111111","100000110110001","100011010011101","100111000001111","100110100110101","100110011101100","000000101011010","100100000011110","000100101101110","000010011101011","000111000100010","000110010010111","100000110010011","000100001000110","100101000010001","000101000001110","100100111010010","100010010100010","000000001000011","000011010111100","000111001000100","000110011001110","100000110100100","100011010001101","100111001010100","000000110110000","100100000010110","000100110100010","100100011101100","100010011001101","000000000101110","000011001001000","100000000100010","100011001111100","100111001000001","000000101100101","000010111101110","000000000000011","000011111100011","100100110000111","100010011000111","000000000101111","100011111000101","000100101000011","100100111111100","100010010101100","000000000010011","000011000101001","000111010110110","000110011001110","000110011010100","000110011011110","100000101101000","000100001100010","100100110101010","000100100101001","100100101010111","100010100001000","000000001010000","000011001000000","000111011000110","000110010011000","100000111100001","000100000111101","100100111110001","000100111000101","000010011101001","100000000001001","100011001111100","000000010000101","000011001001110","000111001011010","000110010010000","000110010011000","100000110111111","100010111110111","100111001111111","000000101101100","000011001001001","000111010010100","100000111101110","000100000101000","100100111101111","100010011010101","100000001110110","100011111011101","100010010011111","100111010010010","100110010111000","000000110100100","100011110110100","000100110100001","100100101010110","100010011010100","100000000101001","000011001100011","000111001011001","100000101100000","100011001101010","100000000110110","000011001011100","000111010110011","100000110110100","000011111010101","000010100001100","000000000000110","000011111101000","100100111001001","000100100111001","000010011010110","000111001010001","000110011100001","000110001101110","000110100100010","100000101111010","000011110011010","100100101010101","000100101110011","000010011100000","000111001110100","000110010010011","100001001010010","100011001000011","100000000010110","000011000111111","000000000011011","100011010010011","000000000101011","000011001110000","000111000100110","000110100000010","100000101111010","100011000010101","100000000111001","100100000111001","000100110101101","000010011110111","000000000110101","100011001100101","100111001110101","100110010100010","100110001001101","000000111010010","000011001101011","000111001000001","000110011101101","000110010101101","100000110001010","100011000110011","100111000101010","000000110111111","100011110100110","100010001010100","100111011100001","000000100100110","000011000101010","000110111100101","100000110110000","000011111101010","100100110001001","100010010111010","100111010010010","000000101100100","000011010011001","100000000011000","100011010111111","000000000000000","000011001110011","100000000011010","100011000111011","000000000001110","100100000001101","100010011001111","000000000011101","000011001001001","000111000100010","000110011000010","100000110010001","000100000100000","100100110011011","000100101111011","000010011110011","000111001011111","100000101100101","100011001101100","100111001100110","000000110010011","100100000111011","100010100001000","100111010100100","100110001011001","000000110001100","000011010100011","000111001111101","100000100100001","100011000101010","100111010110101","000000110000100","100011111000110","100010010111010","000000010010010","000011001100011","000111000000001","000110011101001","000110010010001","100000110010110","100011000100000","000000000010011","000011001111001","100000000001100","000011111110110","100100110100000","000100011100100","000010011100110","000000001000000","100011010111010","100111011001000","100110010100100","100110100101110","000000100101100","000011010011001","000111000111100","100000101001000","000011110101100","100100111000001","100010010111101","100111001000010","100110010101110","000000110100101","100100000001110","100010011110010","000000000011111","000011001001101","000111010000001","000110100010011","000110000111011","100000100100100","000011111010111","100100101000100","000100111111110","100100111111000","000100110100101","000010110101101","100000000001101","100011001000110","100111001010000","100110001111010","000000111100000","100100000111101","000100101111101","100100110000011","000100110010101","000010101110000","000111010000010","000110011101001","100000111001111","100011010111011","000000000110011","000011001011001","000111010010000","100000111001111","000100000111010","000010001010111","000000001100101","000100000110110","100100110010010","100010100010111","100000000011001","100011111101111","100010001111110","100111010101001","100110001111000","000001001001100","000011001000110","000000000011110","100011010010000","100111011010101","000000111111000","000011010010011","000111001000101","000110011010100","000110010111101","100000111111000","100011100100001","100111001101001","000000101111011","100100000100101","100010100000011","100000001110101","000011001000100","000111001110000","100000111011110","100011001001001","100000000010001","000011001011111","000111000001001","100000111001011","000100000011010","000010010011001","000111001110000","000110101001100","100000101100110","100011000100011","000000010011000","100011110110011","000100110110011","100100100011011","100010100000111","100000000101100","000011011101001","000111010000011","000110011001010","000110011101010","000110010111011","000110010111001","000110010110011","100000110111101","000011111000010","000010011001000","100000000100101","100011000001001","000000000001111","100011110111101","000100110010000","100100110011110","000100111101011","100100100111010","000100110011011","000010100111010","000111010000101","100000110000001","100010111011000","000000001100011","000011010100001","000111010000000","000110010101001","000110011000101","000110101000010","000110001001001","100000111000010","100011001110010","100111001011100","100110101000000","100110010101010","100110010011101","000000101011100","100100000010000","100010100011011","100110111111101","100110010110100","100110011011101","000000101011101","100011111111001","000101000000110","100100110000111","100010010110101","100111010110100","000000110100100","000011010011000","100000001011001","000100001001001","100100011111001","000100100110100","000010001000110","100000000000100","000100000110001","100100110011110","100010011010111","000000000000000","100100001000100","000100100101111","100100100110011","100010010111001","100111010110011","000000111011111","100100001010100","000100110010001","100100101101001","100010100000011","100111001111101","000000110011011","100011110000001","100010010101111","100000000011001","100100000001110","100010011011110","100111000010001","100110011011111","100110100000000","000000110101001","100100000000110","000100111001100","100100101011011","100010010000110","100111000111100","000000111000010","000011011100001","000111000011011","100000110110000","000011110010010","100100101011110","100010011001011","100111001111001","100110100111100","000000110100101","100100000010000","000100101000001","100100111100100","100010011111110","100000000010000","000010111111011","000111001011010","100000101110001","100011001111110","100111010010011","000000110101101","100011110111000","100010011101001","100000000011110","000011000001001","000111000100111","000110011110100","000110011000101","000110011111110","000110011111000","100000110000001","100011000110100","000000001100010","000011010001011","000111010000001","100000110011100","100011010110110","100000000100000","000011001111011","100000001000111","000100000011110","000010011100001","000000000000110","100011001010010","000000000000001","000011001100100","000111001100101","000110100001000","000110011000110","100001001000100","000011111100000","100100110001100","100010010001110","000000001011001","000011000101001","000000000110001","100011001010110","100000000001101","000011001101000","100000000000001","000100000001001","100100110001010","000100101101110","100100111011101","000100111011000","000010010111110","000000001011011","100011010100010","100000000100110","000011011000010","000000001011011","100011010101001","100111001011001","100110001110101","000000111101111","000011000010011","000111011001111","100000101101110","000100000001110","000010010111110","000111000100111","100000110010011","000011111101111","000010101100010","000000000001100","000011111110100","000010011001011","000111000111110","000110101010010","100000101110000","000100000000100","100100101010000","100010011001110","100000000000110","000011001000010","100000000100111","000100001100111","100100101100111","000100110011111","100100100101011","100010011001011","100111001010011","000000100111101","000011010000101","100000001011101","100011010100110","100111000101000","100110010110110","000000101100001","000011001001100","000111001110111","000110011011011","100001000001000","100011010110100","100111011011001","000000110010100","100100001101111","100010010011111","100111010100111","100110100010100","100110001011000","100110001000000","100110100000001","000000110010111","000011011100101","000111001000011","100000100101010","100011000110001","000000000000011","100100000010110","100010001011111","000000000101110","100100000101000","100010010110011","100000000111000","100011111110110","100010001101001","000000000100010","000011000110101","000000000010110","100011010010011","100110111100011","000000100100101","100100000101010","000100111001011","100100111001110","100010011001011","000000000101010","100011110101110","000100101011101","000010011000001","000111001000111","100000110100000","000100000010111","100100111000001","100010010011000","000000000011011","000011001000111","000000000010001","100011000100110","000000001000000","100011111010100","100010011010001","100000000101000","000011001110100","000111001001000","000110010110111","100000101011101","100011000001000","000000000100110","000011011101011","000111000000011","000110011001110","000110011010010","100000100110001","000100000100000","000010010110111","000000000100011","100011000111100","000000000001011","100100010000011","100010010001010","100000011100010","000011001101101","000111000000001","000110010110101","100000100111111","000011111011110","000010101001000","000111010011000","000110010111100","100000111010100","000011111011111","000010011100101","000110111001100","100000101110001","100011001010100","100111000110001","000001000011110","100100000010100","000100101011010","000010100011001","000000000111001","100011001101111","100111010001100","100110010111100","100110100010101","100110011001000","000000101110000","000011000110001","000000000111110","000100000000001","000010100100100","000111000100000","100000110001010","000011110111100","000010011110100","000000001010100","000100001000010","100101000100010","000100111000101","000010011001101","000111001111100","000110010101001","100001000000100","000100000111001","100100110111010","100010011100010","000000000001010","100011101011011","000101000101110","100100111101111","100010011101011","100111000100110","000000100010011","000011010110110","000111001010001","000110100100111","100000111010010","000011111000100","100100100000011","100010010100110","100000000010100","100100001000010","000100111100001","100100110000011","100010101011111","100000000111010","000011100100110","000111001100101","100001000011011","100011010011111","100000000011011","100011111010011","000100110001111","100100110010011","100010011001101","100111010100100","100110010000000","000000110000001","000011001001000","000000000001100","100011001101010","100111010001000","000000110100001","000011011101111","000000000100011","000011111010101","000010010010100","000111001010110","100000111111111","000100001110110","000010011011010","100000001001011","100011001011110","100000001011101","100011111011010","000100110001101","000010011001111","000111001111101","100000101100010","100011010011010","100111011000101","000000110010010","100100000110101","000100110110101","000010001010100","000111010011110","100000110000101","100011010101110","100111001111010","000000111001111","100011101100010","100010011100011","000000001011001","100100000110111","100010010111111","100000000001101","000011001111100","100000000100000","000011110100011","100100110101011","000100110110110","100100110111010","100010011011000","100111001001100","100110010101001","100110011111100","100110011011110","000000111010001","100011111101010","100010100100100","100111000000010","100110011110100","000000101101100","000011000001010","100000000000111","100011001101101","100000000010100","000011000110000","100000001101011","000100011000011","100100100111000","000100110000010","000010011000101","000111001111101","000110011001100","000110010100111","100000101011101","100011010110000","000000001111110","000010111110100","000111001010001","000110100000101","000110011010100","000110001101011","100000101011101","000100000001010","000010010011000","000000000011010","000100000110000","100100100001100","100010011010010","100111001111001","100110011101101","100110101001001","000000110111011","000010111100001","100000000010001","000011111101110","100100101100010","000100011100110","000010100001000","000111001000100","000110001111001","100000110011010","000100000001111","000010010110001","000111000000111","100000101001011","100011001011001","100000000101101","100011110110001","100010010110101","100111010111000","100110010100100","000000100100101","000011000100001","000000000001001","000100000011010","100100110010101","000100100011100","000010100000001","000111010111000","000110100011000","000110010100111","100000110110011","100011010101000","000000000010000","000011001110110","100000000110001","100011000101010","100111000101111","000000111000100","000011000110101","000111000001111","000110011110111","100000100111011","100011010111001","100000010001111","000011011000011","000111001100010","000110100011001","100000101011001","100011010110101","100111010000010","100110100000010","100110011000001","100110010000001","100110011001001","100110101010100","000000111101001","100011111111111","000100101111011","000010001000100","000111001111110","100000110001001","000100000010101","100100111011111","000100101101010","100100111010100","100010001011001","100111010011011","000000110001100","100100000111001","000100111010100","100100110011010","000100110011110","100100101011100","000100111000101","000010011111111","100000010001010","000100000001110","100100101011011","100010010110110","100111000101011","100110001000011","100110001111011","100110100010101","100110100000010","100110011010100","000000101101111","000011001100001","000000001001111","100011010001000","100111001111000","100110011011011","000000111000101","000011010101001","100000000001001","100011001111010","100111000101001","100110010011101","100110010101101","000001001101101","100011111111101","000100110101111","100100110011111","000100111000001","100100110111011","000100111011010","000010101000011","000000000000101","100011001101010","100000000100100","100100000011110","000100100101011","100100110011101","100010100000101","000000001010001","000011001110000","000000000000011","100011000001011","100000001110010","000011001111011","000111000100001","000110010100011","000110011011101","000110100000110","000110010010110","000110011110000","000110100101011","100000111010000","100011010100110","100111001100111","000000111000010","100011111111111","000100101100100","100100110010010","000100110100111","000010010110000","000111000011101","000110011101000","000110011001101","000110010110101","000110010100011","100000110111010","100011010011110","100000001000011","100011110101110","000100110001001","000010001011100","000111001000110","000110100010001","000110010101001","000110100111111","000110010011010","000110010011100","000110010001001","000110100011000","100000110111111","100011001001011","100111011010001","000000101110100","100011111010101","000100101000110","100100110010110","100010010101001","000000001110011","100011111010110","100010010001111","100000000010110","100100000100101","000100110011101","000010010010010","000111010101111","000110011111111","100000101011011","000100001010001","000010011000101","000111001000001","100000101110111","000100001001010","100100101100010","100010010001111","000000001100001","000011001111001","000000001001101","000011111111111","100100101100110","100010100100111","000000001100011","000010111110011","000111001110011","000110010110110","000110010000001","100000110000011","100011001010000","000000001011011","100011111110111","100010010100111","000000000001111","100011110100000","000100111100010","000010011001101","000000000001000","100010111110011","100111001110101","100110010010101","100110100000101","100110011111110","000000111010001","100011111010110","100010010001000","100111010001111","100110010001010","100110011000001","000000110010110","100011110010010","000100111110110","100101000101011","100010010110101","100000000110111","000011001010011","000111000111101","000110100110110","000110100011101","100000101110101","100011000111000","100111001001000","000000111000101","100011111101111","100010011011000","000000000100000","100100000010100","000100110000000","000010010111011","000111001100000","000110011001101","000110101110000","000110001111101","100000111011111","000100000001111","100100110011100","100010011111100","100111001010001","000000111001010","100100001001010","000100101111111","000010001111001","000111001101011","100000110001110","000100000101100","000010010000110","000000000010011","100011001101111","000000001011010","000011001111010","100000000100010","000011111110001","000010010101010","000111011000011","000110010101011","000110001100100","100000110100110","100011000011100","100111000111011","000000110100100","000011011011010","000111001000000","000110011011101","000110010010100","000110010011001","100000110101111","100011000111100","100110111100001","100110010011001","100110100010010","100110011011010","000000101110101","000011001010011","000111010110010","000110011100101","100000101011001","100011000111111","100111010011001","000000111010101","000011000001110","000111010011010","100000101110010","100011000011111","100111011000010","100110011011001","000000110011010","000011001101100","000111010011111","100000101101100","000100000101010","000010011011000","000111011010010","000110010110111","000110011010011","100000110111110","100011001101010","100111000110111","000000101001010","100011111110011","000100101101010","000010011111111","000110111100111","000110001001110","100000100110000","100011001110000","100111011100101","000000100101100","100100000000101","100010010111000","000000000010101","000011010101011","000000000010101","100011001101011","000000001000011","100011101111010","000100110011011","100100110101001","000100111011100","000010010101011","100000001100000","100011001101101","000000000001111","100011111110110","000100101010001","100100111000000","000100101101101","100100101011011","000100110010001","000010011110110","000111010001101","000110011000000","000110001001100","000110011100100","100000101101100","000011111001111","000010011001011","000111001001001","100000100101011","100011001101000","000000000001101","100100001000011","000100101101001","000010001110100","000000000101111","000100000100111","100100111001111","100010000010001","100111000101010","100110010110010","000001000010101","100100010011111","100010011010010","100111001100111","100110010111111","000000101010110","100011111011101","000100100001010","000010011010011","000111010000010","000110011001010","000110011100100","000110010011011","100000101110110","100011001111110","100000001101011","000011001010010","000111000111110","100000111011011","000100000100000","100100110010110","000100110001001","000010010101001","000111011010010","100000101001101","000011111110011","000010011010010","000000001100001","100010111110010","100111000011110","000000110000100","100100000100101","100010010011100","100000000110111","000011000100001","000111001001111","000110100001010","100000110001111","100011001010110","000000001001000","000011001110101","100000001001001","000100000110110","100100101111010","100010011010010","100000000011010","000011001000011","000111001100100","100000111001101","000011111011110","100100111111001","000100101111000","100100111000110","100010010100111","000000001011110","100011110111100","000100111011101","000010011111000","000111010001001","000110011111101","100000111001000","100011000110000","100000001001101","100011111010111","000100101100011","000010010001101","100000000011101","100011010111010","100111001100101","000000111100001","100100000010000","000100110111001","100100110001111","000100111101000","100100110100011","100010010111001","000000010011111","000011010110000","000111000101001","100000101010001","100011010100010","100111001100101","100110010111010","100110010010100","100110011100110","100110010101001","100110001011010","000000100011110","000011000100000","000000001001101","000011111101100","000010011001010","000000000111011","000100010001111","100100111101101","100010100000111","100111001101011","100110011001100","100110011000101","000000110000101","000011010110101","100000000111010","000100000001101","100100101011001","000100110110001","000010010100100","000000000000111","100011001111010","100111010001101","100110001110101","100110011011001","100110011110010","000000101101000","000011001101110","100000001100000","000011110010101","100100110001101","100010100100000","100000000011001","000011010011000","000111010100010","000110100110000","100000111011010","000100000110111","000010011100001","000000001010001","100011001011000","000000000110100","100011110110110","100010011100111","100111010000100","100110100100010","100110011010010","100110010110101","100110011111100","100110011001000","000000110000010","100100000011011","100010010011010","100111000110001","100110010000010","100110100010011","000000110010000","100011111010101","100010100100000","000000001111100","100011111110000","100010011110000","000000001000010","100011111100111","000100110100000","000010010100000","100000001110010","100011010100100","100000000101001","100011111100010","000100111000001","100100111001100","000100111001111","100100101101110","100010011010100","100000000111101","000011010100000","100000000001000","000011110111110","000010011011101","000000000100001","100011011000101","000000001111000","000010111011011","100000001101001","100011000010111","100111001010001","100110011101000","000000110011010","000011010010101","100000000111000","000100000111100","100100101101100","100010011001111","000000000001100","000011000111101","000111000101110","100000110110010","100011000100011","100111001110101","000000101111100","000011000100110","100000001001001","000100000000001","000010100010000","000000001001111","100011001000010","100000000010100","000011001001110","000111001111110","000110100001001","000110100001011","100001000100010","100011001101001","100000000111110","000011001000111","000000001110000","100011010011000","100000001101101","000011001110001","000111001011110","000110010110001","000110100000101","000110011110001","000110011100101","100000110101011","000100000010110","000010010111001","000000000001100","000100000100101","100100110000011","000100101101110","100100110111100","100010100010000","000000001000000","100100000000001","100010011110111","100111000111010","000000101111000","000011010000011","000000001100010","000100000111100","100100110100011","100010011010100","000000001111101","000011001011011","000111001111001","100000110000100","000100000111011","100100110001011","000100110110001","100100110000100","100010000011110","000000000111000","000011000101101","100000001001110","000011110010111","100100100100010","000100101100100","000010100001101","000111010001000","000110001101001","100000100010110","100011001000010","100110111110000","100110010110110","000000110100101","000011000100100","000111001101000","100000110010000","000011110011101","100100110011010","000100110100100","000010010011110","000000000011010","100011010110100","100111010001011","100110011000101","100110011110011","000000110110100","100100000010111","100010100000101","000000000111100","100011111011001","000100110111110","000010011111001","000000001000001","100011000100110","100111001100100","000000101111100","100100000000111","100010001111100","100000001001101","000011001000001","000111010101001","000110100000011","000110010101100","100000110100110","100011001110000","100000000010001","000010111001000","100000000011011","100011001010010","000000010011110","000011000000111","100000000101001","100011001111111","100111010100011","000000101101101","100100001111100","100010011010100","100111010000111","100110010101010","000000110011101","000011010101011","000111011001111","100000110010001","000011110101111","100100110001001","100010001110010","100111001101100","000000110110010","000011000100111","000111011001000","000110011100110","000110010110001","000110001100000","000110010100000","100000111011100","000011111100000","100100110000011","000100111001111","100100110001111","100010011000111","000000000011000","100011101010100","100010010110111","100111001011101","100110001100110","000000110011111","000011000111010","000000000111100","100011001111101","000000000001101","000011010011111","000000000110100","100011011001110","100000010011000","000011000111000","000111011010001","000110011011100","100000110100011","100011001110000","100111000100011","100110010110111","000000110111000","100100010000111","000100110001110","000010011001110","000111000101110","100000110011011","100011010001101","100111000101110","000000101110100","000011010111010","000111001100011","100000101011111","100010111010010","000000000000100","000011011000111","000111000100000","000110101000010","000110001111110","100000110011101","100011001111011","100111010110000","100110100100001","100110010100010","100110100100110","100110100100011","000000111100010","000011001100110","000111001111110","000110010010010","100000110100110","100011001010010","100111001011011","000001000001101","000011000111101","100000000001001","100011000110000","100111000101000","000000100011001","000011001001101","000111000111010","100000110011010","000100000100001","000010011101001","000000001001001","100011001001001","000000000010100","100011111000010","000100110110101","100100111101111","100010011000101","100000001101011","100011110111000","000100100010001","100100110111101","100010011000110","100111001101000","100110001010010","000000110011101","100100000100111","000100110111111","100100111100111","100010010101001","000000000010000","100100000011001","000100101110001","100100111100110","000100100011111","100100110110101","100010010011010","100111010010100","000001000000000","000011000101100","000111011110001","000110010011111","000110011010011","100000100111100","100011000010110","100111010010111","100110010011100","100110100010100","100110100111011","000000111000100","100100001110000","100010101010111","100000000000011","000011011000000","000000001001110","000011110011111","000010011001111","000000000110011","100011000100111","100111000000001","100110001100110","100110010010101","000000100111101","000011001101000","100000001011001","100011000010110","000000001110000","000010111100100","000111010011100","000110010110110","100000110111000","100011010011111","100111000010100","000000110110010","000011001011110","000111010000001","000110100001110","000110010010100","100000111001101","100011000111001","100110111111111","000000111101010","100100000000111","000100101000011","000010000110101","000111000101010","000110100010101","100000110111101","000100000010010","100100110001011","100010101011011","000000001010001","000011011101001","000111001100011","000110100001101","000110010011011","100000101110010","000100010001001","000010100100001","100000000101101","000011110111101","000010011010000","000111001010111","100000110011101","100011000010100","100111001011000","100110001100001","000000110010110","100100000001000","100010010011001","100111001001010","100110011011010","100110100110011","000000101010001","100011111011000","100010010101001","100111011000101","100110011000101","100110010101010","100110100011000","100110100001101","000000111100110","100100001110001","100010010101111","100111000100111","000000100100101","000011001011101","000111000011010","000110011010010","100000110110100","100011011010001","000000000101000","000011010001101","000111000111110","000110011101110","100000111110000","000011110110000","000010010000010","000111001011111","100000110111011","100010111101010","100000000000100","100011111011011","000100110111110","100100110000001","100010011000000","100111000010101","100110100011000","000001000000011","000011010010010","000111000011011","000110100010100","000110100011001","100000100101011","100011010000001","000000001101010","000011001110111","000111000000111","100000111001011","000100000111100","000010101000000","000111000011001","000110011000101","100000111000100","100010111101100","100000000111010","000011010111100","000111000111101","100000101100111","000011110101010","100100100111000","100010101011011","100111001010001","000000110110100","100100000110101","100010100001011","100111000111110","000000101010110","000011001100100","100000010110110","000011101111001","000010011001001","000000001001000","100011011010001","000000000101011","100011111011111","100010011110010","100111001100111","100110000111110","100110100100111","100110010101101","100110010111111","000000110101110","000011001100110","000111001111000","000110010111100","100001000000111","000011111011010","100100110001010","000100110101010","000010011110011","000111011110110","100001000000100","000100000101100","100100110010000","100010011001111","100000000101100","000011001011110","000111010010010","100000101111101","100011011001110","100111000101011","100110010111100","100110001010010","100110100010100","100110011111011","100110100111110","100110011001100","100110010001100","100110011101011","000000101110111","000011001010011","100000000001010","000100001000010","100100110011000","000100101111010","000010011110101","000111000001110","000110011110011","100000110100110","000100010001010","100100111000011","000100110110101","000010011010100","100000001000101","100011000101101","100000010010000","000010111101000","100000001010100","100011000010001","100111000100110","100110100011101","100110011011000","000000101101001","100011111110000","000101000100001","100100111010010","100010001001110","100000000011110","000011000111100","000111010001101","100000101101011","100011001010100","100000001011111","000011000111001","100000000111000","100011010000111","100111010011001","100110010110001","000000111011011","100100000010000","000100110111101","000010011111101","000000000001000","100011001111000","100000000100011","000011000011011","100000000010001","100011001011100","100000000001100","000011001110100","000000000000010","100011000111010","100111010001111","100110011010100","000000110101001","000011001001110","000000000010010","100011011011001","000000000011101","000011010000100","100000000000000","000011111101001","000010010110000","100000001101110","000100001000110","000010011110101","000111000011111","100000111111001","000011111100111","100100101101101","100010010010110","100111001000011","000000111001011","100011110001110","000100100101011","000010011101011","100000000000011","000011111001111","000010011111011","100000000000000","000100001001101","000010010001001","000111000101111","100000101111101","100011010011111","100111001011110","000000101111111","000011010101101","000000000011100","100011010000000","100111010001111","000000101111111","000011100000001","100000000000011","000011111110010","000010011000000","000000001100010","000011110001111","100100101010001","100010011111011","100111001111000","100110010100000","100110100001001","100110010110001","000000110010100","000011000001011","000000000001100","000100000100101","100100101110000","000100101110100","000010011001011","000111010001110","100000101110111","000011111100110","000010001111010","000000000010001","000100000010100","000010100101101","000111000000001","100000110110000","000100000011100","000010011000110","000111011101001","100000110110001","000011101100110","100100101101010","100010100100111","000000001010101","100011111100101","000100110000011","100100111011001","100010001010100","100111001010010","000000101111001","000011000111001","000111001011010","000110100011110","100000100011101","000100000000001","000010011101000","000111001111011","000110001100010","000110011010101","100000110111001","100011010000010","100111001110000","100110110001000","100110011111100","000000111001010","000011001101110","100000000100001","000011111101001","000010010000110","100000000101101","000011111011010","000010011000000","000000000100110","100011001100111","100000000000101","000011000110000","000000000111111","100011001010111","100111001000001","000000110100111","000011010011010","000000001100001","100011010000010","000000000100011","100011111010100","100010011001101","000000001111011","000011000100111","000111001000110","000110011010001","000110011001110","100000110101000","000011111100000","000010100000010","100000000000011","100011010011010","000000001101110","100011111000100","000100111111010","000010011001011","000000001111100","000100000111011","100101000001110","100010100011110","000000000100101","000011001011110","100000000001001","100011000100000","100110111111000","100110010110011","000000110100001","100011101101110","100010011001101","100111010000011","000000101110011","100100000101111","000100110011110","100100111010001","100010101000101","100111010111001","000000110110101","100011110111001","000100111100111","000010101100010","000111000100000","100000101000001","000100000000101","000010010101110","000111001001010","100000101011111","100011000111100","100111011011011","100110010001010","100110010010111","000000110001010","000011000100110","100000000110001","000011110101111","000010011001001","000111001001101","000110010111000","100000110001011","000011111101100","100101000000111","000100101110010","000010010101010","000110111110111","100000101100000","100011011110010","000000000011011","000011001010011","000111001001110","100000101101111","000011111101100","100100110101000","000100101100001","100100101010000","100010010001100","000000000101100","000011010001000","000111010010101","000110011111001","100000110000000","000100000101000","100100111000111","100010011001010","000000000100011","000011000110111","000000000000000","000011111110011","100100101001001","100010010101110","100111000011111","000000111000001","000011010100111","000111001100000","000110011010100","000110010100100","000110011100101","000110110010011","100000110010011","100011001101001","100111000101110","000000100110100","000011010101111","000111000101111","100000101110100","100011001010100","100000000000100","100100000101110","100010010110001","000000001001000","000011010010010","000111011000000","000110001110010","000110011001110","000110001110101","100000110010010","000100000100011","100100111001011","000100111101100","100100110111000","100010010100100","100111001111100","100110011111101","000000101101001","100100001011101","000100111111100","100101000111000","000100101000110","000010001001100","100000001010110","100011100011011","100111000111111","000000110011100","000011000100011","000111000010010","000110001110111","000110010111010","000110001001001","000110011100111","100000110011111","000011111101001","100100101101111","000100110101111","000010010110110","000111001101000","100000110100010","000011111010111","100100101010001","000100111100111","100100110010100","000100101010111","000010010000000","000000000010000","100011001110111","100111010011011","000000110100010","000011000011001","000111001111100","000110001100101","100001000111000","000011111110010","000010010001101","000000001100011","000100001011000","100100111000001","000100101011010","000010010111110","100000000010100","000100001011001","000010010110110","000111010110100","000110100011100","000110101101111","100000110110010","000011111100001","100100100101101","100010011111100","100111011011011","100110011000111","000000110111001","100100000010111","100010011100011","100111010111110","100110001011101","100110010111111","100110011110000","000000110110011","000011010011100","100000001000011","000100000001110","000010010101101","000000001101010","100011001011100","100000001001000","000011001011111","000000000011101","100010111011110","100111001100011","100110010100111","000000111100111","000011010000111","100000000111000","000011111110101","100100111000100","100010010011111","000000001100011","000011001100100","000111010101010","100000111000110","100011001011100","100111001110001","000001000000011","000011001111001","000111010011000","100000110101111","100011010001111","000000000011001","100100000110101","000100101000001","100100110101101","000101000000001","000010010110011","000111001110100","000110010100110","000110001001000","000110011001100","000110100111010","000110010110111","100000111100100","100011010100110","000000000010111","000011001001011","000111010100110","100000110101011","000011101111000","100100110110110","100010010011110","100111000100011","100110001111001","000000111011010","100011110111010","000101000010100","100100100110110","000100110100100","100100110111000","100010011011110","000000000101101","100011110110001","000100110001001","100100100110111","100010011111011","100000000011110","100100000011001","000100101101110","000010100000101","100000000001100","100010111101110","100111001100110","000001000010010","000010111001001","000111001111101","100000110000111","000100001111101","000010011011101","000000001110011","000100001111010","000010010100100","100000001001101","000100000110111","100100111001110","000100110001111","000010010100111","000000000000110","000100000100110","000010011111010","000000000001000","100011010100011","100000000110110","000011001111001","100000010001101","000011110110011","000010001100111","000111001010001","100000101111010","000100010011001","000010011001100","100000001000101","000011111100010","100100101111011","100010010001010","100111010000100","000000110011001","000011010110011","000000000001110","000100000000101","000010010110111","100000000011000","100011000100001","100000000100010","100100000000011","000100101010110","100100101110010","100010010111100","100111001001001","000000110010111","100100000110000","100010011010010","100111010111001","100110011100010","000001000101111","000011011010010","000000000111000","100011001001010","000000000110101","100011111100110","000100111010101","100100101001011","100010100001110","100000000001100","000011001100100","000111001000010","100000111011001","000100001010010","000010011111000","100000000111010","100011010101010","100111001001010","100110011111001","100110100011010","100110011011100","100110100000011","000000111010000","100011101101010","100010100111010","000000000110110","100011111100100","100010100000011","000000000111110","000011000101100","000110111101100","100000111100010","000100000100101","100100101111111","100010010001011","000000000011111","000011010111000","100000010000001","100011001111010","100000000010111","100100000000011","100010010000111","100000000101011","100011111101111","100010101001000","100111010100001","000000111010110","000010111110101","000000001011011","000011111100000","000010011101110","000111000011010","000110011111101","100000110011001","000100001010001","100100110111101","100010011111100","100111010010111","100110001001100","000000110000100","100100001101000","100010010001111","100111001100100","100110011100011","000000110111011","100011111000110","100010011110110","000000000000111","000011001010010","100000000100101","100011001000111","000000000101110","100100001011000","100010010000100","100111001011100","100110011011100","100110100110011","000000110001000","100100000000100","000100110100000","100100110110101","000100111010101","100100100110100","000100111101010","100100110101000","100010010110111","100111001001100","000000101110001","100100000000000","100010011110010","100111001100001","100110001100100","100110011011000","100110011111100","100110001110011","100110010010100","100110011101110","100110011111100","000000111110100","100011111111101","100010011000000","000000000010110","000011000111101","000000001000110","100010111001110","100111100000111","100110010111111","000000111010110","100100000110011","000100110011111","100100110001110","100010011110011","000000000101101","000011010110101","000111001110100","100000110000001","100011010001001","100111000011101","000000110010011","000011010000010","000000001001100","000011111101100","000010011000000","000111001101100","000110010111110","100000111101011","000100000011111","000010001101111","000111001010010","100000111110100","000100001010100","000010011010010","000000000011111","000011111101110","100100100110010","100010011100110","100111000011011","100110010000010","000000101110111","000011010000010","000111001101110","000110101010101","000110010001100","000110001100110","000110011100000","100000111011000","000011111011001","100100110000100","100010100100000","100111000100000","000000110110100","000011011000010","000111001010010","100000101011110","000011110110111","100100110001010","100010010000100","100111010010000","000000110011111","000011011010000","100000000110010","100011010101110","100111000101001","000000110011000","100100001000111","100010100000110","000000000010110","000011001110110","100000000010110","100011001010111","100111001000001","000000101101010","100100000010100","000100101101010","100100101000010","000100101000110","000010100110101","100000000100100","000011111111111","100100101011011","100010010011101","100000000010110","100011111000110","000100101001101","100100101000000","100010010000001","000000000000001","100011111100101","100010010001101","100111001111011","000000110111100","000011010010010","000111001111110","000110001110000","000110010110111","100001000011001","000011111100111","100100111001100","100010011010011","100111001001101","000000111001111","000011001011101","000111001101000","000110100001110","000110100100000","000110011011010","000110100000100","100000111001000","100010111111111","100000000101010","000011000110100","000000000100010","000011111111011","100101000000000","000100111011111","100100101101100","000101000000100","000010011011111","000111010010100","000110010000010","000110101000101","100000100000000","000011111100111","100100111000110","000100111011010","000010010000011","000000000001001","000011111110111","000010100000010","100000001111111","100011001011110","000000000010000","100100001110010","100010011010111","100111000111101","100110100011111","000000110000110","100011111110011","000100101110111","000010100110010","000111010011000","100000110111111","000100000010101","100100101010000","100010010111100","100111001000010","100110010100011","000000111001001","100100001010101","100010011111000","100000000010110","000010111111110","100000001011010","100011001001111","100111001001111","000000111010101","000011001111110","100000000110001","100011001100111","100000000101110","100011111000111","000100100110111","000010100000100","000111010000110","100000101100111","000011111011010","100100110001100","100010011001111","100000001100001","100011111100000","100010010110000","100000000110000","000011010110110","000110111110100","100000110110100","100011001111111","100111010010100","100110011110111","000000110111000","100100000111000","000100110011110","000010010110001","100000000001000","000100001111101","100100110111100","000100111010010","100100110010111","000100110011011","000010001010001","000000001000010","100011001011100","100000000011100","100011111111101","100010011010011","000000001110110","100100001000111","000100101110101","100100110001000","100010001010100","100111001010101","100110010000100","000000111001010","000011010010100","000000001010011","000100010010100","100100110010000","000100110000110","100100110001101","100010011100000","100111011111100","000000110010010","100011111110101","000100110000001","000010010111110","000000001010000","000100000000101","000010011001010","000111000111011","100000110111101","000011111111001","100100110010001","000100110110010","000010100110110","000111010111110","100000111100111","100010111110100","100000000111111","000011100001100","000111001110011","100000110110110","100011011101001","100000000011001","000011011001010","100000000011010","100011010000011","100111010111011","000000101001101","000011001000000","000111001111101","000110001000111","100000101101110","000011111100000","100100101100101","000100110011001","100100110110110","100010010101100","100111001000101","000001000011100","000011000010010","100000000101101","000011110110000","000010010100111","000111001000101","000110010110000","100000110110111","100011010000111","100000000001111","100011111100100","000100111100001","100100110110001","000101000001111","100100101100001","100010001111101","100000000111111","100100001110110","000100110101110","000010011100011","100000001101110","100011011000110","000000000010110","100011110111100","100010001110100","100000000111011","100011111011000","000100111000001","000010011001010","100000001000100","100011010101101","100111000110110","100110100111001","000000110000110","100011111110110","000100111100000","000010010110101","000111000001100","000110011100011","100000111001000","100010111110011","100000000111000","000011001110001","000111011101010","000110100010001","000110011001011","100000101111010","100010111001010","100111000001011","100110100100010","100110011000000","100110010000111","100110100110000","000000110101100","100100000000100","100010010111010","100000000110100","100100001110110","000100101010100","100100100100000","000100110010001","000010010001111","000111011000101","100000101011110","000011111001000","000010100010010","000111010101110","100000111001011","100011001000011","100000000011000","000011010110111","100000001010001","100011010000000","000000000110101","000011001100001","000000000100101","100010111110101","100000000011011","100100001000110","100010001100111","100111010000010","100110010111000","000000101110011","000011000000000","000111000101001","100000101000100","100011010000001","100111001110000","100110010111001","100110010000000","000000110100011","100100000010000","000100101100010","000010011110010","000110111011111","000110010000000","100000101101001","000100000011100","000010001111010","000000000100010","000100000011110","100100111100110","100010011010001","000000001100111","100100000011111","100010100100100","000000000001010","100100000100100","000100110000010","100100101111111","100010011010000","100111001111111","100110100001111","100110100000001","000000101010111","100100000100111","100010001011010","100111001011100","000000101110110","000011001011110","000000000001111","000100000010001","100100110000100","000100111100000","000010010110110","000000000010110","100011010001110","100111011011110","100110011110001","100110001110000","100110011100011","000000111011011","000011010001101","100000000100110","100010111101010","000000000111000","000011010100000","000111000101011","000110010100010","100000101101111","000100001001101","100100110011011","000101000001000","100100110100001","100010010011110","000000000000000","000011010101101","100000000010101","100011001101000","100000001100001","100011111101100","000100110011111","100100101110111","100010010110110","100000000101011","000011010010001","000000010101001","100011010001111","000000000111100","000011001000000","100000000111010","000011110110111","000010011110010","000000000000010","000100000111000","100100110100101","100010100011000","100000000001100","000011001100001","000111010001110","000110001111110","000110001010101","000110011101010","100000111001011","000011111100000","000010011110000","000111001100111","000110011010111","000110100011001","000110100010001","100000110011001","100011010001000","100111010110011","000000110101110","000011011111100","000111010101010","000110011011011","100000111100000","100011010110101","100111010001000","100110110111111","000000110110100","000011010110110","000000000000111","000011111101010","000010100100100");
  variable Y,ERR,TEMP,TEMP_E : sfixed(7 downto -22);
  variable PERCENT_ERROR,I,N,COUNT: integer; 
  variable ARRAY_COUNT :integer range -1 to 4999 := -1;
  variable STEP_SIZE : sfixed(3 downto -11):= "000000000001010";

    begin
    if rising_edge(CLK) then
         ARRAY_COUNT := ARRAY_COUNT+1;
         if(ARRAY_COUNT = 4999) then
         ARRAY_COUNT := 0;
         end if ; 
        for I in 9 downto 1 loop
            IN_FRAME(I)<= IN_FRAME(I-1);
        end loop;
        IN_FRAME(0) <= INPUT_ARRAY(ARRAY_COUNT);
        
        for N in 9 downto 0 loop 
        Y:= WEIGHTS(N)*IN_FRAME(N);
        end loop ;
        
        OUT_SIG <= Y;
        --TEMP_E := to_sfixed(CORRECT_SIGNAL,7,-22) - Y; 
        ERR := resize(arg => (EXPECTED_ARRAY(n)-IN_FRAME(0)),left_index=>7,right_index=> -22,round_style=>fixed_round,overflow_style=> fixed_wrap);
        
        for I in 9 downto 0 loop
        --TEMP := WEIGHTS(I)+ E*IN_FRAME(I);
        WEIGHTS(I)<= resize(arg => WEIGHTS(I)+ STEP_SIZE*ERR*IN_FRAME(I),left_index=>3,right_index=> -11,round_style=>fixed_round,overflow_style=> fixed_wrap); -- ADD STEP SIZE HERE
        end loop;
        
        PERCENT_ERROR := to_integer(ERR*100);
        
        if(PERCENT_ERROR < 1) then
            COUNT := COUNT + 1;
            else
            COUNT := 0;
        end if;
        
        if(COUNT = 100) then 
            LED_LOW_ERROR <= '1' ;
            else
            LED_LOW_ERROR <= '0' ;
        end if;
    end if ;
end process;
end EQUALIZER;
